`include "../Common/scoreboard_base.sv"


module scramble_descramble_top;

    /* Parameters */
    localparam DATA_WIDTH = 32;
    localparam SCRAMBLER = 0;
    localparam DESCRAMBLER = 1;

    /* Signal Descriptions */
    logic clk;
    logic i_reset_n;

    // Scrambler Interface 
    logic i_rx_data_valid;
    logic [DATA_WIDTH-1:0] i_rx_data;
    logic o_tx_trdy;
    logic o_tx_data_valid;
    logic [DATA_WIDTH-1:0] o_tx_data;
    logic i_rx_trdy;

    // De-scrambler Interface
    logic i_rx_data_valid_grbx;
    logic [DATA_WIDTH-1:0] i_rx_data_grbx;
    logic o_tx_trdy_dscrmbl;
    logic o_tx_data_valid_dscrmbl;
    logic [DATA_WIDTH-1:0] o_tx_data_dscrmbl;
    logic i_rx_trdy_dcoder;    

    /* Queue Declarations */
    logic [31:0] tx_queue[$];

    /* Scoreboard Declaration */
    scoreboard_base scb = new();

    /* DUT Instantiation */
    scrambler #(
        .DATA_WIDTH(DATA_WIDTH),
        .DESCRAMBLE(SCRAMBLER) // Set to descramble
    ) Scrambler_DUT (
        .i_clk(clk),
        .i_reset_n(i_reset_n),

        // Encoder-to-Scrambler Interface
        .i_rx_data(i_rx_data),
        .i_rx_data_valid(i_rx_data_valid),
        .o_tx_trdy(o_tx_trdy),

        // Scrambler-to-Gearbox Interface
        .o_tx_data(o_tx_data),
        .o_tx_data_valid(o_tx_data_valid),
        .i_rx_trdy(i_rx_trdy)
    );

    scrambler #(
        .DATA_WIDTH(DATA_WIDTH),
        .DESCRAMBLE(DESCRAMBLER) // Set to descramble
    ) Descrambler_DUT (
        .i_clk(clk),
        .i_reset_n(i_reset_n),

        // Gearbox to Scrambler
        .i_rx_data(i_rx_data_grbx),
        .i_rx_data_valid(i_rx_data_valid_grbx),
        .o_tx_trdy(o_tx_trdy_dscrmbl),

        // Scrambler to decoder
        .o_tx_data(o_tx_data_dscrmbl),
        .o_tx_data_valid(o_tx_data_valid_dscrmbl),
        .i_rx_trdy(i_rx_trdy_dcoder)
    );    

    // Loopback Logic
    assign i_rx_data_grbx = o_tx_data;
    assign i_rx_data_valid_grbx = o_tx_data_valid;

    /* Clock Instantiation */

    always #10 clk = ~clk;

    initial begin
        clk = 1'b0;
    end

    /* Generate and transmit data to the scrambler */
    task generate_data();
        logic [31:0] data_in;
        
        data_in = $urandom;
        i_rx_data_valid <= 1'b1;
        i_rx_data <= data_in; 
        tx_queue.push_back(data_in);
        //$display("Data Pushed into queue: %0h", data_in);
        @(posedge clk); 
    endtask : generate_data

    // Grab the input data generated and validate this with the expected data 
    // generated by the golden model
    function validate_data();
        logic [31:0] input_data;
        logic [57:0] lfsr_golden = {58{1'b1}};

        if (o_tx_data_valid_dscrmbl & i_rx_trdy_dcoder) begin
            // Grab data from queue
            input_data = tx_queue.pop_front();
            //$display("Data sampled from queue: %0h", input_data);

            assert(o_tx_data_dscrmbl == input_data) begin
                $display("PASSED: Input = 0x%08h, Output = 0x%08h", input_data, o_tx_data);
                scb.record_success();
            end else begin
                $display("FAILED: Input = 0x%08h, Output = 0x%08h", input_data, o_tx_data);     
                scb.record_failure();           
            end
        end
    endfunction: validate_data

    /* Stimulus/Test */
    initial begin
        i_rx_data_valid = 1'b0;
        i_rx_data = 32'h0;
        i_rx_trdy = 1'b1;
        i_rx_trdy_dcoder = 1'b1;
        i_rx_data_grbx = 32'b0;
        i_rx_data_valid_grbx = 1'b0;


        // Initial Reset for design
        i_reset_n = 1'b0; #10;
        @(posedge clk)
        i_reset_n = 1'b1;        

        fork
            begin
                for(int i = 0; i < $urandom_range(200, 500); i++) begin                    
                    generate_data();
                end
                i_rx_data_valid <= 1'b0;
                @(posedge clk);
            end
            begin
                while(1) begin
                    validate_data();                     
                    @(posedge clk);
                end
            end
        join_any

        scb.print_summary();

        #100;
        $finish;

    end


endmodule : scramble_descramble_top
