`include "../Common/scoreboard_base.sv"


module descrambler_top;

    /* Parameters */
    localparam DATA_WIDTH = 32;
    localparam SCRAMBLER_BYPASS = 0;

    /* Signal Descriptions */
    logic clk;
    logic i_reset_n;

    logic i_rx_data_valid;
    logic [DATA_WIDTH-1:0] i_rx_data;
    logic o_tx_trdy;
    logic o_tx_data_valid;
    logic [DATA_WIDTH-1:0] o_tx_data;
    logic i_rx_trdy;

    /* Queue Declarations */
    logic [31:0] tx_queue[$];

    /* Scoreboard Declaration */
    scoreboard_base scb = new();

    /* DUT Instantiation */
    scrambler #(
        .DATA_WIDTH(DATA_WIDTH),
        .DESCRAMBLE(1) // Set to descramble
    ) DUT (
        .i_clk(clk),
        .i_reset_n(i_reset_n),

        // Encoder-to-Scrambler Interface
        .i_rx_data(i_rx_data),
        .i_rx_data_valid(i_rx_data_valid),
        .o_tx_trdy(o_tx_trdy),

        // Scrambler-to-Gearbox Interface
        .o_tx_data(o_tx_data),
        .o_tx_data_valid(o_tx_data_valid),
        .i_rx_trdy(i_rx_trdy)
    );

    /* Clock Instantiation */

    always #10 clk = ~clk;

    initial begin
        clk = 1'b0;
    end

    /* Golden Model */
    function automatic [31:0] scramble_golden_model (
        input  logic [31:0] data_in,
        inout  logic [57:0] lfsr
    );
        logic [31:0] data_out;
        logic feedback;
        int i;

        for (i = 0; i < 32; i++) begin
            // Shift LFSR and insert new feedback bit
            lfsr = {lfsr[56:0], data_in[i]};            
            // Scramble input bit using MSB of LFSR
            data_out[i] = data_in[i] ^ lfsr[57] ^ lfsr[38];
        end

        return data_out;

    endfunction    

    /* Generate and transmit data to the scrambler */
    task generate_data();
        logic [31:0] data_in;
        
        data_in = $urandom;
        i_rx_data_valid <= 1'b1;
        i_rx_data <= data_in; 
        tx_queue.push_back(data_in);
        @(posedge clk); 
    endtask : generate_data

    // Grab the input data generated and validate this with the expected data 
    // generated by the golden model
    function validate_data();
        logic [31:0] expected_out, input_data;
        logic [57:0] lfsr_golden = {58{1'b1}};

        if (o_tx_data_valid & i_rx_trdy) begin
            // Grab data from queue
            input_data = tx_queue.pop_front();
            // Generate expected data
            expected_out = scramble_golden_model(input_data, lfsr_golden);

            assert(o_tx_data == expected_out) begin
                $display("PASSED: Input = 0x%08h, Output = 0x%08h", input_data, o_tx_data);
                scb.record_success();
            end else begin
                $display("FAILED: Input = 0x%08h, Output = 0x%08h, Expected: %0h", input_data, o_tx_data, expected_out);     
                scb.record_failure();           
            end
        end
    endfunction: validate_data

    task scrambler_test_case();
        fork
            begin
                for(int i = 0; i < $urandom_range(50, 100); i++) begin                    
                    generate_data();
                end
                i_rx_data_valid <= 1'b0;
                @(posedge clk);
            end
            begin
                while(1) begin
                    validate_data();                     
                    @(posedge clk);
                end
            end
        join_any
    endtask : scrambler_test_case

    /* Stimulus/Test */
    initial begin
        i_rx_data_valid = 1'b0;
        i_rx_data = 32'h0;
        i_rx_trdy = 1'b1;

        // Initial Reset for design
        i_reset_n = 1'b0; #10;
        @(posedge clk)
        i_reset_n = 1'b1;        

        fork
            begin
                for(int i = 0; i < $urandom_range(50, 100); i++) begin                    
                    generate_data();
                end
                i_rx_data_valid <= 1'b0;
                @(posedge clk);
            end
            begin
                while(1) begin
                    validate_data();                     
                    @(posedge clk);
                end
            end
        join_any

        scb.print_summary();

        #100;
        $finish;

    end


endmodule : descrambler_top