
package decoder_pkg;


endpackage : decoder_pkg